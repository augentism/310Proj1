library verilog;
use verilog.vl_types.all;
entity muxor16 is
    port(
        y               : out    vl_logic_vector(15 downto 0);
        a               : in     vl_logic_vector(15 downto 0);
        b               : in     vl_logic_vector(15 downto 0)
    );
end muxor16;
